-- Nios_System_A1.vhd

-- Generated using ACDS version 18.1 625

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity Nios_System_A1 is
	port (
		button_pio_external_connection_export    : in    std_logic_vector(3 downto 0)  := (others => '0'); --    button_pio_external_connection.export
		clocks_ref_clk_clk                       : in    std_logic                     := '0';             --                    clocks_ref_clk.clk
		clocks_ref_reset_reset                   : in    std_logic                     := '0';             --                  clocks_ref_reset.reset
		clocks_sdram_clk_clk                     : out   std_logic;                                        --                  clocks_sdram_clk.clk
		led_pio_external_connection_export       : out   std_logic_vector(7 downto 0);                     --       led_pio_external_connection.export
		sdram_wire_addr                          : out   std_logic_vector(12 downto 0);                    --                        sdram_wire.addr
		sdram_wire_ba                            : out   std_logic_vector(1 downto 0);                     --                                  .ba
		sdram_wire_cas_n                         : out   std_logic;                                        --                                  .cas_n
		sdram_wire_cke                           : out   std_logic;                                        --                                  .cke
		sdram_wire_cs_n                          : out   std_logic;                                        --                                  .cs_n
		sdram_wire_dq                            : inout std_logic_vector(15 downto 0) := (others => '0'); --                                  .dq
		sdram_wire_dqm                           : out   std_logic_vector(1 downto 0);                     --                                  .dqm
		sdram_wire_ras_n                         : out   std_logic;                                        --                                  .ras_n
		sdram_wire_we_n                          : out   std_logic;                                        --                                  .we_n
		segment_1_pio_external_connection_export : out   std_logic_vector(6 downto 0);                     -- segment_1_pio_external_connection.export
		segment_2_pio_external_connection_export : out   std_logic_vector(6 downto 0);                     -- segment_2_pio_external_connection.export
		segment_3_pio_external_connection_export : out   std_logic_vector(6 downto 0);                     -- segment_3_pio_external_connection.export
		segment_4_pio_external_connection_export : out   std_logic_vector(6 downto 0);                     -- segment_4_pio_external_connection.export
		switch_pio_external_connection_export    : in    std_logic_vector(7 downto 0)  := (others => '0')  --    switch_pio_external_connection.export
	);
end entity Nios_System_A1;

architecture rtl of Nios_System_A1 is
	component Nios_System_A1_BUTTON_pio is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			in_port    : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- export
			irq        : out std_logic                                         -- irq
		);
	end component Nios_System_A1_BUTTON_pio;

	component Nios_System_A1_LED_pio is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(7 downto 0)                      -- export
		);
	end component Nios_System_A1_LED_pio;

	component SIMD_MULTI_Instruction is
		port (
			dataa  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- dataa
			datab  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- datab
			result : out std_logic_vector(31 downto 0)                     -- result
		);
	end component SIMD_MULTI_Instruction;

	component Nios_System_A1_Segment_1 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(6 downto 0)                      -- export
		);
	end component Nios_System_A1_Segment_1;

	component Nios_System_A1_Switches_0_7 is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic_vector(7 downto 0)  := (others => 'X')  -- export
		);
	end component Nios_System_A1_Switches_0_7;

	component Nios_System_A1_clocks is
		port (
			ref_clk_clk        : in  std_logic := 'X'; -- clk
			ref_reset_reset    : in  std_logic := 'X'; -- reset
			sys_clk_clk        : out std_logic;        -- clk
			sdram_clk_clk      : out std_logic;        -- clk
			reset_source_reset : out std_logic         -- reset
		);
	end component Nios_System_A1_clocks;

	component Nios_System_A1_cpu is
		port (
			clk                                 : in  std_logic                     := 'X';             -- clk
			reset_n                             : in  std_logic                     := 'X';             -- reset_n
			reset_req                           : in  std_logic                     := 'X';             -- reset_req
			d_address                           : out std_logic_vector(27 downto 0);                    -- address
			d_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                              : out std_logic;                                        -- read
			d_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			d_write                             : out std_logic;                                        -- write
			d_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			debug_mem_slave_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                           : out std_logic_vector(27 downto 0);                    -- address
			i_read                              : out std_logic;                                        -- read
			i_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			debug_reset_request                 : out std_logic;                                        -- reset
			debug_mem_slave_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			debug_mem_slave_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			debug_mem_slave_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			debug_mem_slave_read                : in  std_logic                     := 'X';             -- read
			debug_mem_slave_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			debug_mem_slave_waitrequest         : out std_logic;                                        -- waitrequest
			debug_mem_slave_write               : in  std_logic                     := 'X';             -- write
			debug_mem_slave_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			E_ci_combo_result                   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- result
			E_ci_combo_a                        : out std_logic_vector(4 downto 0);                     -- a
			E_ci_combo_b                        : out std_logic_vector(4 downto 0);                     -- b
			E_ci_combo_c                        : out std_logic_vector(4 downto 0);                     -- c
			E_ci_combo_dataa                    : out std_logic_vector(31 downto 0);                    -- dataa
			E_ci_combo_datab                    : out std_logic_vector(31 downto 0);                    -- datab
			E_ci_combo_estatus                  : out std_logic;                                        -- estatus
			E_ci_combo_ipending                 : out std_logic_vector(31 downto 0);                    -- ipending
			E_ci_combo_n                        : out std_logic_vector(7 downto 0);                     -- n
			E_ci_combo_readra                   : out std_logic;                                        -- readra
			E_ci_combo_readrb                   : out std_logic;                                        -- readrb
			E_ci_combo_writerc                  : out std_logic                                         -- writerc
		);
	end component Nios_System_A1_cpu;

	component Nios_System_A1_high_res_timer is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			writedata  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata   : out std_logic_vector(15 downto 0);                    -- readdata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write_n    : in  std_logic                     := 'X';             -- write_n
			irq        : out std_logic                                         -- irq
		);
	end component Nios_System_A1_high_res_timer;

	component Nios_System_A1_jtag_uart is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component Nios_System_A1_jtag_uart;

	component Nios_System_A1_onchip_memory is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			address    : in  std_logic_vector(12 downto 0) := (others => 'X'); -- address
			clken      : in  std_logic                     := 'X';             -- clken
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write      : in  std_logic                     := 'X';             -- write
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset      : in  std_logic                     := 'X';             -- reset
			reset_req  : in  std_logic                     := 'X';             -- reset_req
			freeze     : in  std_logic                     := 'X'              -- freeze
		);
	end component Nios_System_A1_onchip_memory;

	component Nios_System_A1_sdram is
		port (
			clk            : in    std_logic                     := 'X';             -- clk
			reset_n        : in    std_logic                     := 'X';             -- reset_n
			az_addr        : in    std_logic_vector(24 downto 0) := (others => 'X'); -- address
			az_be_n        : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- byteenable_n
			az_cs          : in    std_logic                     := 'X';             -- chipselect
			az_data        : in    std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			az_rd_n        : in    std_logic                     := 'X';             -- read_n
			az_wr_n        : in    std_logic                     := 'X';             -- write_n
			za_data        : out   std_logic_vector(15 downto 0);                    -- readdata
			za_valid       : out   std_logic;                                        -- readdatavalid
			za_waitrequest : out   std_logic;                                        -- waitrequest
			zs_addr        : out   std_logic_vector(12 downto 0);                    -- export
			zs_ba          : out   std_logic_vector(1 downto 0);                     -- export
			zs_cas_n       : out   std_logic;                                        -- export
			zs_cke         : out   std_logic;                                        -- export
			zs_cs_n        : out   std_logic;                                        -- export
			zs_dq          : inout std_logic_vector(15 downto 0) := (others => 'X'); -- export
			zs_dqm         : out   std_logic_vector(1 downto 0);                     -- export
			zs_ras_n       : out   std_logic;                                        -- export
			zs_we_n        : out   std_logic                                         -- export
		);
	end component Nios_System_A1_sdram;

	component altera_customins_master_translator is
		generic (
			SHARED_COMB_AND_MULTI : integer := 0
		);
		port (
			ci_slave_dataa            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- dataa
			ci_slave_datab            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- datab
			ci_slave_result           : out std_logic_vector(31 downto 0);                    -- result
			ci_slave_n                : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- n
			ci_slave_readra           : in  std_logic                     := 'X';             -- readra
			ci_slave_readrb           : in  std_logic                     := 'X';             -- readrb
			ci_slave_writerc          : in  std_logic                     := 'X';             -- writerc
			ci_slave_a                : in  std_logic_vector(4 downto 0)  := (others => 'X'); -- a
			ci_slave_b                : in  std_logic_vector(4 downto 0)  := (others => 'X'); -- b
			ci_slave_c                : in  std_logic_vector(4 downto 0)  := (others => 'X'); -- c
			ci_slave_ipending         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- ipending
			ci_slave_estatus          : in  std_logic                     := 'X';             -- estatus
			comb_ci_master_dataa      : out std_logic_vector(31 downto 0);                    -- dataa
			comb_ci_master_datab      : out std_logic_vector(31 downto 0);                    -- datab
			comb_ci_master_result     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- result
			comb_ci_master_n          : out std_logic_vector(7 downto 0);                     -- n
			comb_ci_master_readra     : out std_logic;                                        -- readra
			comb_ci_master_readrb     : out std_logic;                                        -- readrb
			comb_ci_master_writerc    : out std_logic;                                        -- writerc
			comb_ci_master_a          : out std_logic_vector(4 downto 0);                     -- a
			comb_ci_master_b          : out std_logic_vector(4 downto 0);                     -- b
			comb_ci_master_c          : out std_logic_vector(4 downto 0);                     -- c
			comb_ci_master_ipending   : out std_logic_vector(31 downto 0);                    -- ipending
			comb_ci_master_estatus    : out std_logic;                                        -- estatus
			ci_slave_multi_clk        : in  std_logic                     := 'X';             -- clk
			ci_slave_multi_reset      : in  std_logic                     := 'X';             -- reset
			ci_slave_multi_clken      : in  std_logic                     := 'X';             -- clk_en
			ci_slave_multi_reset_req  : in  std_logic                     := 'X';             -- reset_req
			ci_slave_multi_start      : in  std_logic                     := 'X';             -- start
			ci_slave_multi_done       : out std_logic;                                        -- done
			ci_slave_multi_dataa      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- multi_dataa
			ci_slave_multi_datab      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- multi_datab
			ci_slave_multi_result     : out std_logic_vector(31 downto 0);                    -- multi_result
			ci_slave_multi_n          : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- multi_n
			ci_slave_multi_readra     : in  std_logic                     := 'X';             -- multi_readra
			ci_slave_multi_readrb     : in  std_logic                     := 'X';             -- multi_readrb
			ci_slave_multi_writerc    : in  std_logic                     := 'X';             -- multi_writerc
			ci_slave_multi_a          : in  std_logic_vector(4 downto 0)  := (others => 'X'); -- multi_a
			ci_slave_multi_b          : in  std_logic_vector(4 downto 0)  := (others => 'X'); -- multi_b
			ci_slave_multi_c          : in  std_logic_vector(4 downto 0)  := (others => 'X'); -- multi_c
			multi_ci_master_clk       : out std_logic;                                        -- clk
			multi_ci_master_reset     : out std_logic;                                        -- reset
			multi_ci_master_clken     : out std_logic;                                        -- clk_en
			multi_ci_master_reset_req : out std_logic;                                        -- reset_req
			multi_ci_master_start     : out std_logic;                                        -- start
			multi_ci_master_done      : in  std_logic                     := 'X';             -- done
			multi_ci_master_dataa     : out std_logic_vector(31 downto 0);                    -- dataa
			multi_ci_master_datab     : out std_logic_vector(31 downto 0);                    -- datab
			multi_ci_master_result    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- result
			multi_ci_master_n         : out std_logic_vector(7 downto 0);                     -- n
			multi_ci_master_readra    : out std_logic;                                        -- readra
			multi_ci_master_readrb    : out std_logic;                                        -- readrb
			multi_ci_master_writerc   : out std_logic;                                        -- writerc
			multi_ci_master_a         : out std_logic_vector(4 downto 0);                     -- a
			multi_ci_master_b         : out std_logic_vector(4 downto 0);                     -- b
			multi_ci_master_c         : out std_logic_vector(4 downto 0)                      -- c
		);
	end component altera_customins_master_translator;

	component Nios_System_A1_cpu_custom_instruction_master_comb_xconnect is
		port (
			ci_slave_dataa      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- dataa
			ci_slave_datab      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- datab
			ci_slave_result     : out std_logic_vector(31 downto 0);                    -- result
			ci_slave_n          : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- n
			ci_slave_readra     : in  std_logic                     := 'X';             -- readra
			ci_slave_readrb     : in  std_logic                     := 'X';             -- readrb
			ci_slave_writerc    : in  std_logic                     := 'X';             -- writerc
			ci_slave_a          : in  std_logic_vector(4 downto 0)  := (others => 'X'); -- a
			ci_slave_b          : in  std_logic_vector(4 downto 0)  := (others => 'X'); -- b
			ci_slave_c          : in  std_logic_vector(4 downto 0)  := (others => 'X'); -- c
			ci_slave_ipending   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- ipending
			ci_slave_estatus    : in  std_logic                     := 'X';             -- estatus
			ci_master0_dataa    : out std_logic_vector(31 downto 0);                    -- dataa
			ci_master0_datab    : out std_logic_vector(31 downto 0);                    -- datab
			ci_master0_result   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- result
			ci_master0_n        : out std_logic_vector(7 downto 0);                     -- n
			ci_master0_readra   : out std_logic;                                        -- readra
			ci_master0_readrb   : out std_logic;                                        -- readrb
			ci_master0_writerc  : out std_logic;                                        -- writerc
			ci_master0_a        : out std_logic_vector(4 downto 0);                     -- a
			ci_master0_b        : out std_logic_vector(4 downto 0);                     -- b
			ci_master0_c        : out std_logic_vector(4 downto 0);                     -- c
			ci_master0_ipending : out std_logic_vector(31 downto 0);                    -- ipending
			ci_master0_estatus  : out std_logic                                         -- estatus
		);
	end component Nios_System_A1_cpu_custom_instruction_master_comb_xconnect;

	component altera_customins_slave_translator is
		generic (
			N_WIDTH          : integer := 8;
			USE_DONE         : integer := 1;
			NUM_FIXED_CYCLES : integer := 2
		);
		port (
			ci_slave_dataa      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- dataa
			ci_slave_datab      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- datab
			ci_slave_result     : out std_logic_vector(31 downto 0);                    -- result
			ci_slave_n          : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- n
			ci_slave_readra     : in  std_logic                     := 'X';             -- readra
			ci_slave_readrb     : in  std_logic                     := 'X';             -- readrb
			ci_slave_writerc    : in  std_logic                     := 'X';             -- writerc
			ci_slave_a          : in  std_logic_vector(4 downto 0)  := (others => 'X'); -- a
			ci_slave_b          : in  std_logic_vector(4 downto 0)  := (others => 'X'); -- b
			ci_slave_c          : in  std_logic_vector(4 downto 0)  := (others => 'X'); -- c
			ci_slave_ipending   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- ipending
			ci_slave_estatus    : in  std_logic                     := 'X';             -- estatus
			ci_master_dataa     : out std_logic_vector(31 downto 0);                    -- dataa
			ci_master_datab     : out std_logic_vector(31 downto 0);                    -- datab
			ci_master_result    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- result
			ci_master_n         : out std_logic_vector(7 downto 0);                     -- n
			ci_master_readra    : out std_logic;                                        -- readra
			ci_master_readrb    : out std_logic;                                        -- readrb
			ci_master_writerc   : out std_logic;                                        -- writerc
			ci_master_a         : out std_logic_vector(4 downto 0);                     -- a
			ci_master_b         : out std_logic_vector(4 downto 0);                     -- b
			ci_master_c         : out std_logic_vector(4 downto 0);                     -- c
			ci_master_ipending  : out std_logic_vector(31 downto 0);                    -- ipending
			ci_master_estatus   : out std_logic;                                        -- estatus
			ci_master_clk       : out std_logic;                                        -- clk
			ci_master_clken     : out std_logic;                                        -- clk_en
			ci_master_reset_req : out std_logic;                                        -- reset_req
			ci_master_reset     : out std_logic;                                        -- reset
			ci_master_start     : out std_logic;                                        -- start
			ci_master_done      : in  std_logic                     := 'X';             -- done
			ci_slave_clk        : in  std_logic                     := 'X';             -- clk
			ci_slave_clken      : in  std_logic                     := 'X';             -- clk_en
			ci_slave_reset_req  : in  std_logic                     := 'X';             -- reset_req
			ci_slave_reset      : in  std_logic                     := 'X';             -- reset
			ci_slave_start      : in  std_logic                     := 'X';             -- start
			ci_slave_done       : out std_logic                                         -- done
		);
	end component altera_customins_slave_translator;

	component Nios_System_A1_mm_interconnect_0 is
		port (
			clocks_sys_clk_clk                      : in  std_logic                     := 'X';             -- clk
			cpu_reset_reset_bridge_in_reset_reset   : in  std_logic                     := 'X';             -- reset
			cpu_data_master_address                 : in  std_logic_vector(27 downto 0) := (others => 'X'); -- address
			cpu_data_master_waitrequest             : out std_logic;                                        -- waitrequest
			cpu_data_master_byteenable              : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			cpu_data_master_read                    : in  std_logic                     := 'X';             -- read
			cpu_data_master_readdata                : out std_logic_vector(31 downto 0);                    -- readdata
			cpu_data_master_write                   : in  std_logic                     := 'X';             -- write
			cpu_data_master_writedata               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			cpu_data_master_debugaccess             : in  std_logic                     := 'X';             -- debugaccess
			cpu_instruction_master_address          : in  std_logic_vector(27 downto 0) := (others => 'X'); -- address
			cpu_instruction_master_waitrequest      : out std_logic;                                        -- waitrequest
			cpu_instruction_master_read             : in  std_logic                     := 'X';             -- read
			cpu_instruction_master_readdata         : out std_logic_vector(31 downto 0);                    -- readdata
			BUTTON_pio_s1_address                   : out std_logic_vector(1 downto 0);                     -- address
			BUTTON_pio_s1_write                     : out std_logic;                                        -- write
			BUTTON_pio_s1_readdata                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			BUTTON_pio_s1_writedata                 : out std_logic_vector(31 downto 0);                    -- writedata
			BUTTON_pio_s1_chipselect                : out std_logic;                                        -- chipselect
			cpu_debug_mem_slave_address             : out std_logic_vector(8 downto 0);                     -- address
			cpu_debug_mem_slave_write               : out std_logic;                                        -- write
			cpu_debug_mem_slave_read                : out std_logic;                                        -- read
			cpu_debug_mem_slave_readdata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			cpu_debug_mem_slave_writedata           : out std_logic_vector(31 downto 0);                    -- writedata
			cpu_debug_mem_slave_byteenable          : out std_logic_vector(3 downto 0);                     -- byteenable
			cpu_debug_mem_slave_waitrequest         : in  std_logic                     := 'X';             -- waitrequest
			cpu_debug_mem_slave_debugaccess         : out std_logic;                                        -- debugaccess
			high_res_timer_s1_address               : out std_logic_vector(2 downto 0);                     -- address
			high_res_timer_s1_write                 : out std_logic;                                        -- write
			high_res_timer_s1_readdata              : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			high_res_timer_s1_writedata             : out std_logic_vector(15 downto 0);                    -- writedata
			high_res_timer_s1_chipselect            : out std_logic;                                        -- chipselect
			jtag_uart_avalon_jtag_slave_address     : out std_logic_vector(0 downto 0);                     -- address
			jtag_uart_avalon_jtag_slave_write       : out std_logic;                                        -- write
			jtag_uart_avalon_jtag_slave_read        : out std_logic;                                        -- read
			jtag_uart_avalon_jtag_slave_readdata    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			jtag_uart_avalon_jtag_slave_writedata   : out std_logic_vector(31 downto 0);                    -- writedata
			jtag_uart_avalon_jtag_slave_waitrequest : in  std_logic                     := 'X';             -- waitrequest
			jtag_uart_avalon_jtag_slave_chipselect  : out std_logic;                                        -- chipselect
			LED_pio_s1_address                      : out std_logic_vector(1 downto 0);                     -- address
			LED_pio_s1_write                        : out std_logic;                                        -- write
			LED_pio_s1_readdata                     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			LED_pio_s1_writedata                    : out std_logic_vector(31 downto 0);                    -- writedata
			LED_pio_s1_chipselect                   : out std_logic;                                        -- chipselect
			onchip_memory_s1_address                : out std_logic_vector(12 downto 0);                    -- address
			onchip_memory_s1_write                  : out std_logic;                                        -- write
			onchip_memory_s1_readdata               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			onchip_memory_s1_writedata              : out std_logic_vector(31 downto 0);                    -- writedata
			onchip_memory_s1_byteenable             : out std_logic_vector(3 downto 0);                     -- byteenable
			onchip_memory_s1_chipselect             : out std_logic;                                        -- chipselect
			onchip_memory_s1_clken                  : out std_logic;                                        -- clken
			sdram_s1_address                        : out std_logic_vector(24 downto 0);                    -- address
			sdram_s1_write                          : out std_logic;                                        -- write
			sdram_s1_read                           : out std_logic;                                        -- read
			sdram_s1_readdata                       : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			sdram_s1_writedata                      : out std_logic_vector(15 downto 0);                    -- writedata
			sdram_s1_byteenable                     : out std_logic_vector(1 downto 0);                     -- byteenable
			sdram_s1_readdatavalid                  : in  std_logic                     := 'X';             -- readdatavalid
			sdram_s1_waitrequest                    : in  std_logic                     := 'X';             -- waitrequest
			sdram_s1_chipselect                     : out std_logic;                                        -- chipselect
			Segment_1_s1_address                    : out std_logic_vector(1 downto 0);                     -- address
			Segment_1_s1_write                      : out std_logic;                                        -- write
			Segment_1_s1_readdata                   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			Segment_1_s1_writedata                  : out std_logic_vector(31 downto 0);                    -- writedata
			Segment_1_s1_chipselect                 : out std_logic;                                        -- chipselect
			Segment_2_s1_address                    : out std_logic_vector(1 downto 0);                     -- address
			Segment_2_s1_write                      : out std_logic;                                        -- write
			Segment_2_s1_readdata                   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			Segment_2_s1_writedata                  : out std_logic_vector(31 downto 0);                    -- writedata
			Segment_2_s1_chipselect                 : out std_logic;                                        -- chipselect
			Segment_3_s1_address                    : out std_logic_vector(1 downto 0);                     -- address
			Segment_3_s1_write                      : out std_logic;                                        -- write
			Segment_3_s1_readdata                   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			Segment_3_s1_writedata                  : out std_logic_vector(31 downto 0);                    -- writedata
			Segment_3_s1_chipselect                 : out std_logic;                                        -- chipselect
			Segment_4_s1_address                    : out std_logic_vector(1 downto 0);                     -- address
			Segment_4_s1_write                      : out std_logic;                                        -- write
			Segment_4_s1_readdata                   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			Segment_4_s1_writedata                  : out std_logic_vector(31 downto 0);                    -- writedata
			Segment_4_s1_chipselect                 : out std_logic;                                        -- chipselect
			Switches_0_7_s1_address                 : out std_logic_vector(1 downto 0);                     -- address
			Switches_0_7_s1_readdata                : in  std_logic_vector(31 downto 0) := (others => 'X')  -- readdata
		);
	end component Nios_System_A1_mm_interconnect_0;

	component Nios_System_A1_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			receiver1_irq : in  std_logic                     := 'X'; -- irq
			receiver2_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component Nios_System_A1_irq_mapper;

	component altera_reset_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_in1      : in  std_logic := 'X'; -- reset
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component altera_reset_controller;

	signal clocks_sys_clk_clk                                                    : std_logic;                     -- clocks:sys_clk_clk -> [BUTTON_pio:clk, LED_pio:clk, Segment_1:clk, Segment_2:clk, Segment_3:clk, Segment_4:clk, Switches_0_7:clk, cpu:clk, high_res_timer:clk, irq_mapper:clk, jtag_uart:clk, mm_interconnect_0:clocks_sys_clk_clk, onchip_memory:clk, rst_controller:clk, sdram:clk]
	signal cpu_custom_instruction_master_result                                  : std_logic_vector(31 downto 0); -- cpu_custom_instruction_master_translator:ci_slave_result -> cpu:E_ci_combo_result
	signal cpu_custom_instruction_master_readra                                  : std_logic;                     -- cpu:E_ci_combo_readra -> cpu_custom_instruction_master_translator:ci_slave_readra
	signal cpu_custom_instruction_master_a                                       : std_logic_vector(4 downto 0);  -- cpu:E_ci_combo_a -> cpu_custom_instruction_master_translator:ci_slave_a
	signal cpu_custom_instruction_master_b                                       : std_logic_vector(4 downto 0);  -- cpu:E_ci_combo_b -> cpu_custom_instruction_master_translator:ci_slave_b
	signal cpu_custom_instruction_master_c                                       : std_logic_vector(4 downto 0);  -- cpu:E_ci_combo_c -> cpu_custom_instruction_master_translator:ci_slave_c
	signal cpu_custom_instruction_master_readrb                                  : std_logic;                     -- cpu:E_ci_combo_readrb -> cpu_custom_instruction_master_translator:ci_slave_readrb
	signal cpu_custom_instruction_master_estatus                                 : std_logic;                     -- cpu:E_ci_combo_estatus -> cpu_custom_instruction_master_translator:ci_slave_estatus
	signal cpu_custom_instruction_master_ipending                                : std_logic_vector(31 downto 0); -- cpu:E_ci_combo_ipending -> cpu_custom_instruction_master_translator:ci_slave_ipending
	signal cpu_custom_instruction_master_datab                                   : std_logic_vector(31 downto 0); -- cpu:E_ci_combo_datab -> cpu_custom_instruction_master_translator:ci_slave_datab
	signal cpu_custom_instruction_master_dataa                                   : std_logic_vector(31 downto 0); -- cpu:E_ci_combo_dataa -> cpu_custom_instruction_master_translator:ci_slave_dataa
	signal cpu_custom_instruction_master_writerc                                 : std_logic;                     -- cpu:E_ci_combo_writerc -> cpu_custom_instruction_master_translator:ci_slave_writerc
	signal cpu_custom_instruction_master_n                                       : std_logic_vector(7 downto 0);  -- cpu:E_ci_combo_n -> cpu_custom_instruction_master_translator:ci_slave_n
	signal cpu_custom_instruction_master_translator_comb_ci_master_result        : std_logic_vector(31 downto 0); -- cpu_custom_instruction_master_comb_xconnect:ci_slave_result -> cpu_custom_instruction_master_translator:comb_ci_master_result
	signal cpu_custom_instruction_master_translator_comb_ci_master_readra        : std_logic;                     -- cpu_custom_instruction_master_translator:comb_ci_master_readra -> cpu_custom_instruction_master_comb_xconnect:ci_slave_readra
	signal cpu_custom_instruction_master_translator_comb_ci_master_a             : std_logic_vector(4 downto 0);  -- cpu_custom_instruction_master_translator:comb_ci_master_a -> cpu_custom_instruction_master_comb_xconnect:ci_slave_a
	signal cpu_custom_instruction_master_translator_comb_ci_master_b             : std_logic_vector(4 downto 0);  -- cpu_custom_instruction_master_translator:comb_ci_master_b -> cpu_custom_instruction_master_comb_xconnect:ci_slave_b
	signal cpu_custom_instruction_master_translator_comb_ci_master_readrb        : std_logic;                     -- cpu_custom_instruction_master_translator:comb_ci_master_readrb -> cpu_custom_instruction_master_comb_xconnect:ci_slave_readrb
	signal cpu_custom_instruction_master_translator_comb_ci_master_c             : std_logic_vector(4 downto 0);  -- cpu_custom_instruction_master_translator:comb_ci_master_c -> cpu_custom_instruction_master_comb_xconnect:ci_slave_c
	signal cpu_custom_instruction_master_translator_comb_ci_master_estatus       : std_logic;                     -- cpu_custom_instruction_master_translator:comb_ci_master_estatus -> cpu_custom_instruction_master_comb_xconnect:ci_slave_estatus
	signal cpu_custom_instruction_master_translator_comb_ci_master_ipending      : std_logic_vector(31 downto 0); -- cpu_custom_instruction_master_translator:comb_ci_master_ipending -> cpu_custom_instruction_master_comb_xconnect:ci_slave_ipending
	signal cpu_custom_instruction_master_translator_comb_ci_master_datab         : std_logic_vector(31 downto 0); -- cpu_custom_instruction_master_translator:comb_ci_master_datab -> cpu_custom_instruction_master_comb_xconnect:ci_slave_datab
	signal cpu_custom_instruction_master_translator_comb_ci_master_dataa         : std_logic_vector(31 downto 0); -- cpu_custom_instruction_master_translator:comb_ci_master_dataa -> cpu_custom_instruction_master_comb_xconnect:ci_slave_dataa
	signal cpu_custom_instruction_master_translator_comb_ci_master_writerc       : std_logic;                     -- cpu_custom_instruction_master_translator:comb_ci_master_writerc -> cpu_custom_instruction_master_comb_xconnect:ci_slave_writerc
	signal cpu_custom_instruction_master_translator_comb_ci_master_n             : std_logic_vector(7 downto 0);  -- cpu_custom_instruction_master_translator:comb_ci_master_n -> cpu_custom_instruction_master_comb_xconnect:ci_slave_n
	signal cpu_custom_instruction_master_comb_xconnect_ci_master0_result         : std_logic_vector(31 downto 0); -- cpu_custom_instruction_master_comb_slave_translator0:ci_slave_result -> cpu_custom_instruction_master_comb_xconnect:ci_master0_result
	signal cpu_custom_instruction_master_comb_xconnect_ci_master0_readra         : std_logic;                     -- cpu_custom_instruction_master_comb_xconnect:ci_master0_readra -> cpu_custom_instruction_master_comb_slave_translator0:ci_slave_readra
	signal cpu_custom_instruction_master_comb_xconnect_ci_master0_a              : std_logic_vector(4 downto 0);  -- cpu_custom_instruction_master_comb_xconnect:ci_master0_a -> cpu_custom_instruction_master_comb_slave_translator0:ci_slave_a
	signal cpu_custom_instruction_master_comb_xconnect_ci_master0_b              : std_logic_vector(4 downto 0);  -- cpu_custom_instruction_master_comb_xconnect:ci_master0_b -> cpu_custom_instruction_master_comb_slave_translator0:ci_slave_b
	signal cpu_custom_instruction_master_comb_xconnect_ci_master0_readrb         : std_logic;                     -- cpu_custom_instruction_master_comb_xconnect:ci_master0_readrb -> cpu_custom_instruction_master_comb_slave_translator0:ci_slave_readrb
	signal cpu_custom_instruction_master_comb_xconnect_ci_master0_c              : std_logic_vector(4 downto 0);  -- cpu_custom_instruction_master_comb_xconnect:ci_master0_c -> cpu_custom_instruction_master_comb_slave_translator0:ci_slave_c
	signal cpu_custom_instruction_master_comb_xconnect_ci_master0_estatus        : std_logic;                     -- cpu_custom_instruction_master_comb_xconnect:ci_master0_estatus -> cpu_custom_instruction_master_comb_slave_translator0:ci_slave_estatus
	signal cpu_custom_instruction_master_comb_xconnect_ci_master0_ipending       : std_logic_vector(31 downto 0); -- cpu_custom_instruction_master_comb_xconnect:ci_master0_ipending -> cpu_custom_instruction_master_comb_slave_translator0:ci_slave_ipending
	signal cpu_custom_instruction_master_comb_xconnect_ci_master0_datab          : std_logic_vector(31 downto 0); -- cpu_custom_instruction_master_comb_xconnect:ci_master0_datab -> cpu_custom_instruction_master_comb_slave_translator0:ci_slave_datab
	signal cpu_custom_instruction_master_comb_xconnect_ci_master0_dataa          : std_logic_vector(31 downto 0); -- cpu_custom_instruction_master_comb_xconnect:ci_master0_dataa -> cpu_custom_instruction_master_comb_slave_translator0:ci_slave_dataa
	signal cpu_custom_instruction_master_comb_xconnect_ci_master0_writerc        : std_logic;                     -- cpu_custom_instruction_master_comb_xconnect:ci_master0_writerc -> cpu_custom_instruction_master_comb_slave_translator0:ci_slave_writerc
	signal cpu_custom_instruction_master_comb_xconnect_ci_master0_n              : std_logic_vector(7 downto 0);  -- cpu_custom_instruction_master_comb_xconnect:ci_master0_n -> cpu_custom_instruction_master_comb_slave_translator0:ci_slave_n
	signal cpu_custom_instruction_master_comb_slave_translator0_ci_master_result : std_logic_vector(31 downto 0); -- SIMD_MULTI_0:result -> cpu_custom_instruction_master_comb_slave_translator0:ci_master_result
	signal cpu_custom_instruction_master_comb_slave_translator0_ci_master_datab  : std_logic_vector(31 downto 0); -- cpu_custom_instruction_master_comb_slave_translator0:ci_master_datab -> SIMD_MULTI_0:datab
	signal cpu_custom_instruction_master_comb_slave_translator0_ci_master_dataa  : std_logic_vector(31 downto 0); -- cpu_custom_instruction_master_comb_slave_translator0:ci_master_dataa -> SIMD_MULTI_0:dataa
	signal cpu_data_master_readdata                                              : std_logic_vector(31 downto 0); -- mm_interconnect_0:cpu_data_master_readdata -> cpu:d_readdata
	signal cpu_data_master_waitrequest                                           : std_logic;                     -- mm_interconnect_0:cpu_data_master_waitrequest -> cpu:d_waitrequest
	signal cpu_data_master_debugaccess                                           : std_logic;                     -- cpu:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:cpu_data_master_debugaccess
	signal cpu_data_master_address                                               : std_logic_vector(27 downto 0); -- cpu:d_address -> mm_interconnect_0:cpu_data_master_address
	signal cpu_data_master_byteenable                                            : std_logic_vector(3 downto 0);  -- cpu:d_byteenable -> mm_interconnect_0:cpu_data_master_byteenable
	signal cpu_data_master_read                                                  : std_logic;                     -- cpu:d_read -> mm_interconnect_0:cpu_data_master_read
	signal cpu_data_master_write                                                 : std_logic;                     -- cpu:d_write -> mm_interconnect_0:cpu_data_master_write
	signal cpu_data_master_writedata                                             : std_logic_vector(31 downto 0); -- cpu:d_writedata -> mm_interconnect_0:cpu_data_master_writedata
	signal cpu_instruction_master_readdata                                       : std_logic_vector(31 downto 0); -- mm_interconnect_0:cpu_instruction_master_readdata -> cpu:i_readdata
	signal cpu_instruction_master_waitrequest                                    : std_logic;                     -- mm_interconnect_0:cpu_instruction_master_waitrequest -> cpu:i_waitrequest
	signal cpu_instruction_master_address                                        : std_logic_vector(27 downto 0); -- cpu:i_address -> mm_interconnect_0:cpu_instruction_master_address
	signal cpu_instruction_master_read                                           : std_logic;                     -- cpu:i_read -> mm_interconnect_0:cpu_instruction_master_read
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect              : std_logic;                     -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata                : std_logic_vector(31 downto 0); -- jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest             : std_logic;                     -- jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_address                 : std_logic_vector(0 downto 0);  -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_read                    : std_logic;                     -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> mm_interconnect_0_jtag_uart_avalon_jtag_slave_read:in
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_write                   : std_logic;                     -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> mm_interconnect_0_jtag_uart_avalon_jtag_slave_write:in
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata               : std_logic_vector(31 downto 0); -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	signal mm_interconnect_0_cpu_debug_mem_slave_readdata                        : std_logic_vector(31 downto 0); -- cpu:debug_mem_slave_readdata -> mm_interconnect_0:cpu_debug_mem_slave_readdata
	signal mm_interconnect_0_cpu_debug_mem_slave_waitrequest                     : std_logic;                     -- cpu:debug_mem_slave_waitrequest -> mm_interconnect_0:cpu_debug_mem_slave_waitrequest
	signal mm_interconnect_0_cpu_debug_mem_slave_debugaccess                     : std_logic;                     -- mm_interconnect_0:cpu_debug_mem_slave_debugaccess -> cpu:debug_mem_slave_debugaccess
	signal mm_interconnect_0_cpu_debug_mem_slave_address                         : std_logic_vector(8 downto 0);  -- mm_interconnect_0:cpu_debug_mem_slave_address -> cpu:debug_mem_slave_address
	signal mm_interconnect_0_cpu_debug_mem_slave_read                            : std_logic;                     -- mm_interconnect_0:cpu_debug_mem_slave_read -> cpu:debug_mem_slave_read
	signal mm_interconnect_0_cpu_debug_mem_slave_byteenable                      : std_logic_vector(3 downto 0);  -- mm_interconnect_0:cpu_debug_mem_slave_byteenable -> cpu:debug_mem_slave_byteenable
	signal mm_interconnect_0_cpu_debug_mem_slave_write                           : std_logic;                     -- mm_interconnect_0:cpu_debug_mem_slave_write -> cpu:debug_mem_slave_write
	signal mm_interconnect_0_cpu_debug_mem_slave_writedata                       : std_logic_vector(31 downto 0); -- mm_interconnect_0:cpu_debug_mem_slave_writedata -> cpu:debug_mem_slave_writedata
	signal mm_interconnect_0_onchip_memory_s1_chipselect                         : std_logic;                     -- mm_interconnect_0:onchip_memory_s1_chipselect -> onchip_memory:chipselect
	signal mm_interconnect_0_onchip_memory_s1_readdata                           : std_logic_vector(31 downto 0); -- onchip_memory:readdata -> mm_interconnect_0:onchip_memory_s1_readdata
	signal mm_interconnect_0_onchip_memory_s1_address                            : std_logic_vector(12 downto 0); -- mm_interconnect_0:onchip_memory_s1_address -> onchip_memory:address
	signal mm_interconnect_0_onchip_memory_s1_byteenable                         : std_logic_vector(3 downto 0);  -- mm_interconnect_0:onchip_memory_s1_byteenable -> onchip_memory:byteenable
	signal mm_interconnect_0_onchip_memory_s1_write                              : std_logic;                     -- mm_interconnect_0:onchip_memory_s1_write -> onchip_memory:write
	signal mm_interconnect_0_onchip_memory_s1_writedata                          : std_logic_vector(31 downto 0); -- mm_interconnect_0:onchip_memory_s1_writedata -> onchip_memory:writedata
	signal mm_interconnect_0_onchip_memory_s1_clken                              : std_logic;                     -- mm_interconnect_0:onchip_memory_s1_clken -> onchip_memory:clken
	signal mm_interconnect_0_led_pio_s1_chipselect                               : std_logic;                     -- mm_interconnect_0:LED_pio_s1_chipselect -> LED_pio:chipselect
	signal mm_interconnect_0_led_pio_s1_readdata                                 : std_logic_vector(31 downto 0); -- LED_pio:readdata -> mm_interconnect_0:LED_pio_s1_readdata
	signal mm_interconnect_0_led_pio_s1_address                                  : std_logic_vector(1 downto 0);  -- mm_interconnect_0:LED_pio_s1_address -> LED_pio:address
	signal mm_interconnect_0_led_pio_s1_write                                    : std_logic;                     -- mm_interconnect_0:LED_pio_s1_write -> mm_interconnect_0_led_pio_s1_write:in
	signal mm_interconnect_0_led_pio_s1_writedata                                : std_logic_vector(31 downto 0); -- mm_interconnect_0:LED_pio_s1_writedata -> LED_pio:writedata
	signal mm_interconnect_0_sdram_s1_chipselect                                 : std_logic;                     -- mm_interconnect_0:sdram_s1_chipselect -> sdram:az_cs
	signal mm_interconnect_0_sdram_s1_readdata                                   : std_logic_vector(15 downto 0); -- sdram:za_data -> mm_interconnect_0:sdram_s1_readdata
	signal mm_interconnect_0_sdram_s1_waitrequest                                : std_logic;                     -- sdram:za_waitrequest -> mm_interconnect_0:sdram_s1_waitrequest
	signal mm_interconnect_0_sdram_s1_address                                    : std_logic_vector(24 downto 0); -- mm_interconnect_0:sdram_s1_address -> sdram:az_addr
	signal mm_interconnect_0_sdram_s1_read                                       : std_logic;                     -- mm_interconnect_0:sdram_s1_read -> mm_interconnect_0_sdram_s1_read:in
	signal mm_interconnect_0_sdram_s1_byteenable                                 : std_logic_vector(1 downto 0);  -- mm_interconnect_0:sdram_s1_byteenable -> mm_interconnect_0_sdram_s1_byteenable:in
	signal mm_interconnect_0_sdram_s1_readdatavalid                              : std_logic;                     -- sdram:za_valid -> mm_interconnect_0:sdram_s1_readdatavalid
	signal mm_interconnect_0_sdram_s1_write                                      : std_logic;                     -- mm_interconnect_0:sdram_s1_write -> mm_interconnect_0_sdram_s1_write:in
	signal mm_interconnect_0_sdram_s1_writedata                                  : std_logic_vector(15 downto 0); -- mm_interconnect_0:sdram_s1_writedata -> sdram:az_data
	signal mm_interconnect_0_high_res_timer_s1_chipselect                        : std_logic;                     -- mm_interconnect_0:high_res_timer_s1_chipselect -> high_res_timer:chipselect
	signal mm_interconnect_0_high_res_timer_s1_readdata                          : std_logic_vector(15 downto 0); -- high_res_timer:readdata -> mm_interconnect_0:high_res_timer_s1_readdata
	signal mm_interconnect_0_high_res_timer_s1_address                           : std_logic_vector(2 downto 0);  -- mm_interconnect_0:high_res_timer_s1_address -> high_res_timer:address
	signal mm_interconnect_0_high_res_timer_s1_write                             : std_logic;                     -- mm_interconnect_0:high_res_timer_s1_write -> mm_interconnect_0_high_res_timer_s1_write:in
	signal mm_interconnect_0_high_res_timer_s1_writedata                         : std_logic_vector(15 downto 0); -- mm_interconnect_0:high_res_timer_s1_writedata -> high_res_timer:writedata
	signal mm_interconnect_0_button_pio_s1_chipselect                            : std_logic;                     -- mm_interconnect_0:BUTTON_pio_s1_chipselect -> BUTTON_pio:chipselect
	signal mm_interconnect_0_button_pio_s1_readdata                              : std_logic_vector(31 downto 0); -- BUTTON_pio:readdata -> mm_interconnect_0:BUTTON_pio_s1_readdata
	signal mm_interconnect_0_button_pio_s1_address                               : std_logic_vector(1 downto 0);  -- mm_interconnect_0:BUTTON_pio_s1_address -> BUTTON_pio:address
	signal mm_interconnect_0_button_pio_s1_write                                 : std_logic;                     -- mm_interconnect_0:BUTTON_pio_s1_write -> mm_interconnect_0_button_pio_s1_write:in
	signal mm_interconnect_0_button_pio_s1_writedata                             : std_logic_vector(31 downto 0); -- mm_interconnect_0:BUTTON_pio_s1_writedata -> BUTTON_pio:writedata
	signal mm_interconnect_0_switches_0_7_s1_readdata                            : std_logic_vector(31 downto 0); -- Switches_0_7:readdata -> mm_interconnect_0:Switches_0_7_s1_readdata
	signal mm_interconnect_0_switches_0_7_s1_address                             : std_logic_vector(1 downto 0);  -- mm_interconnect_0:Switches_0_7_s1_address -> Switches_0_7:address
	signal mm_interconnect_0_segment_1_s1_chipselect                             : std_logic;                     -- mm_interconnect_0:Segment_1_s1_chipselect -> Segment_1:chipselect
	signal mm_interconnect_0_segment_1_s1_readdata                               : std_logic_vector(31 downto 0); -- Segment_1:readdata -> mm_interconnect_0:Segment_1_s1_readdata
	signal mm_interconnect_0_segment_1_s1_address                                : std_logic_vector(1 downto 0);  -- mm_interconnect_0:Segment_1_s1_address -> Segment_1:address
	signal mm_interconnect_0_segment_1_s1_write                                  : std_logic;                     -- mm_interconnect_0:Segment_1_s1_write -> mm_interconnect_0_segment_1_s1_write:in
	signal mm_interconnect_0_segment_1_s1_writedata                              : std_logic_vector(31 downto 0); -- mm_interconnect_0:Segment_1_s1_writedata -> Segment_1:writedata
	signal mm_interconnect_0_segment_2_s1_chipselect                             : std_logic;                     -- mm_interconnect_0:Segment_2_s1_chipselect -> Segment_2:chipselect
	signal mm_interconnect_0_segment_2_s1_readdata                               : std_logic_vector(31 downto 0); -- Segment_2:readdata -> mm_interconnect_0:Segment_2_s1_readdata
	signal mm_interconnect_0_segment_2_s1_address                                : std_logic_vector(1 downto 0);  -- mm_interconnect_0:Segment_2_s1_address -> Segment_2:address
	signal mm_interconnect_0_segment_2_s1_write                                  : std_logic;                     -- mm_interconnect_0:Segment_2_s1_write -> mm_interconnect_0_segment_2_s1_write:in
	signal mm_interconnect_0_segment_2_s1_writedata                              : std_logic_vector(31 downto 0); -- mm_interconnect_0:Segment_2_s1_writedata -> Segment_2:writedata
	signal mm_interconnect_0_segment_3_s1_chipselect                             : std_logic;                     -- mm_interconnect_0:Segment_3_s1_chipselect -> Segment_3:chipselect
	signal mm_interconnect_0_segment_3_s1_readdata                               : std_logic_vector(31 downto 0); -- Segment_3:readdata -> mm_interconnect_0:Segment_3_s1_readdata
	signal mm_interconnect_0_segment_3_s1_address                                : std_logic_vector(1 downto 0);  -- mm_interconnect_0:Segment_3_s1_address -> Segment_3:address
	signal mm_interconnect_0_segment_3_s1_write                                  : std_logic;                     -- mm_interconnect_0:Segment_3_s1_write -> mm_interconnect_0_segment_3_s1_write:in
	signal mm_interconnect_0_segment_3_s1_writedata                              : std_logic_vector(31 downto 0); -- mm_interconnect_0:Segment_3_s1_writedata -> Segment_3:writedata
	signal mm_interconnect_0_segment_4_s1_chipselect                             : std_logic;                     -- mm_interconnect_0:Segment_4_s1_chipselect -> Segment_4:chipselect
	signal mm_interconnect_0_segment_4_s1_readdata                               : std_logic_vector(31 downto 0); -- Segment_4:readdata -> mm_interconnect_0:Segment_4_s1_readdata
	signal mm_interconnect_0_segment_4_s1_address                                : std_logic_vector(1 downto 0);  -- mm_interconnect_0:Segment_4_s1_address -> Segment_4:address
	signal mm_interconnect_0_segment_4_s1_write                                  : std_logic;                     -- mm_interconnect_0:Segment_4_s1_write -> mm_interconnect_0_segment_4_s1_write:in
	signal mm_interconnect_0_segment_4_s1_writedata                              : std_logic_vector(31 downto 0); -- mm_interconnect_0:Segment_4_s1_writedata -> Segment_4:writedata
	signal irq_mapper_receiver0_irq                                              : std_logic;                     -- jtag_uart:av_irq -> irq_mapper:receiver0_irq
	signal irq_mapper_receiver1_irq                                              : std_logic;                     -- high_res_timer:irq -> irq_mapper:receiver1_irq
	signal irq_mapper_receiver2_irq                                              : std_logic;                     -- BUTTON_pio:irq -> irq_mapper:receiver2_irq
	signal cpu_irq_irq                                                           : std_logic_vector(31 downto 0); -- irq_mapper:sender_irq -> cpu:irq
	signal rst_controller_reset_out_reset                                        : std_logic;                     -- rst_controller:reset_out -> [irq_mapper:reset, mm_interconnect_0:cpu_reset_reset_bridge_in_reset_reset, onchip_memory:reset, rst_controller_reset_out_reset:in, rst_translator:in_reset]
	signal rst_controller_reset_out_reset_req                                    : std_logic;                     -- rst_controller:reset_req -> [cpu:reset_req, onchip_memory:reset_req, rst_translator:reset_req_in]
	signal cpu_debug_reset_request_reset                                         : std_logic;                     -- cpu:debug_reset_request -> rst_controller:reset_in0
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv          : std_logic;                     -- mm_interconnect_0_jtag_uart_avalon_jtag_slave_read:inv -> jtag_uart:av_read_n
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv         : std_logic;                     -- mm_interconnect_0_jtag_uart_avalon_jtag_slave_write:inv -> jtag_uart:av_write_n
	signal mm_interconnect_0_led_pio_s1_write_ports_inv                          : std_logic;                     -- mm_interconnect_0_led_pio_s1_write:inv -> LED_pio:write_n
	signal mm_interconnect_0_sdram_s1_read_ports_inv                             : std_logic;                     -- mm_interconnect_0_sdram_s1_read:inv -> sdram:az_rd_n
	signal mm_interconnect_0_sdram_s1_byteenable_ports_inv                       : std_logic_vector(1 downto 0);  -- mm_interconnect_0_sdram_s1_byteenable:inv -> sdram:az_be_n
	signal mm_interconnect_0_sdram_s1_write_ports_inv                            : std_logic;                     -- mm_interconnect_0_sdram_s1_write:inv -> sdram:az_wr_n
	signal mm_interconnect_0_high_res_timer_s1_write_ports_inv                   : std_logic;                     -- mm_interconnect_0_high_res_timer_s1_write:inv -> high_res_timer:write_n
	signal mm_interconnect_0_button_pio_s1_write_ports_inv                       : std_logic;                     -- mm_interconnect_0_button_pio_s1_write:inv -> BUTTON_pio:write_n
	signal mm_interconnect_0_segment_1_s1_write_ports_inv                        : std_logic;                     -- mm_interconnect_0_segment_1_s1_write:inv -> Segment_1:write_n
	signal mm_interconnect_0_segment_2_s1_write_ports_inv                        : std_logic;                     -- mm_interconnect_0_segment_2_s1_write:inv -> Segment_2:write_n
	signal mm_interconnect_0_segment_3_s1_write_ports_inv                        : std_logic;                     -- mm_interconnect_0_segment_3_s1_write:inv -> Segment_3:write_n
	signal mm_interconnect_0_segment_4_s1_write_ports_inv                        : std_logic;                     -- mm_interconnect_0_segment_4_s1_write:inv -> Segment_4:write_n
	signal rst_controller_reset_out_reset_ports_inv                              : std_logic;                     -- rst_controller_reset_out_reset:inv -> [BUTTON_pio:reset_n, LED_pio:reset_n, Segment_1:reset_n, Segment_2:reset_n, Segment_3:reset_n, Segment_4:reset_n, Switches_0_7:reset_n, cpu:reset_n, high_res_timer:reset_n, jtag_uart:rst_n, sdram:reset_n]

begin

	button_pio : component Nios_System_A1_BUTTON_pio
		port map (
			clk        => clocks_sys_clk_clk,                              --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,        --               reset.reset_n
			address    => mm_interconnect_0_button_pio_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_button_pio_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_button_pio_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_button_pio_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_button_pio_s1_readdata,        --                    .readdata
			in_port    => button_pio_external_connection_export,           -- external_connection.export
			irq        => irq_mapper_receiver2_irq                         --                 irq.irq
		);

	led_pio : component Nios_System_A1_LED_pio
		port map (
			clk        => clocks_sys_clk_clk,                           --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,     --               reset.reset_n
			address    => mm_interconnect_0_led_pio_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_led_pio_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_led_pio_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_led_pio_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_led_pio_s1_readdata,        --                    .readdata
			out_port   => led_pio_external_connection_export            -- external_connection.export
		);

	simd_multi_0 : component SIMD_MULTI_Instruction
		port map (
			dataa  => cpu_custom_instruction_master_comb_slave_translator0_ci_master_dataa,  -- nios_custom_instruction_slave.dataa
			datab  => cpu_custom_instruction_master_comb_slave_translator0_ci_master_datab,  --                              .datab
			result => cpu_custom_instruction_master_comb_slave_translator0_ci_master_result  --                              .result
		);

	segment_1 : component Nios_System_A1_Segment_1
		port map (
			clk        => clocks_sys_clk_clk,                             --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,       --               reset.reset_n
			address    => mm_interconnect_0_segment_1_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_segment_1_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_segment_1_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_segment_1_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_segment_1_s1_readdata,        --                    .readdata
			out_port   => segment_1_pio_external_connection_export        -- external_connection.export
		);

	segment_2 : component Nios_System_A1_Segment_1
		port map (
			clk        => clocks_sys_clk_clk,                             --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,       --               reset.reset_n
			address    => mm_interconnect_0_segment_2_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_segment_2_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_segment_2_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_segment_2_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_segment_2_s1_readdata,        --                    .readdata
			out_port   => segment_2_pio_external_connection_export        -- external_connection.export
		);

	segment_3 : component Nios_System_A1_Segment_1
		port map (
			clk        => clocks_sys_clk_clk,                             --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,       --               reset.reset_n
			address    => mm_interconnect_0_segment_3_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_segment_3_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_segment_3_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_segment_3_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_segment_3_s1_readdata,        --                    .readdata
			out_port   => segment_3_pio_external_connection_export        -- external_connection.export
		);

	segment_4 : component Nios_System_A1_Segment_1
		port map (
			clk        => clocks_sys_clk_clk,                             --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,       --               reset.reset_n
			address    => mm_interconnect_0_segment_4_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_segment_4_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_segment_4_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_segment_4_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_segment_4_s1_readdata,        --                    .readdata
			out_port   => segment_4_pio_external_connection_export        -- external_connection.export
		);

	switches_0_7 : component Nios_System_A1_Switches_0_7
		port map (
			clk      => clocks_sys_clk_clk,                         --                 clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,   --               reset.reset_n
			address  => mm_interconnect_0_switches_0_7_s1_address,  --                  s1.address
			readdata => mm_interconnect_0_switches_0_7_s1_readdata, --                    .readdata
			in_port  => switch_pio_external_connection_export       -- external_connection.export
		);

	clocks : component Nios_System_A1_clocks
		port map (
			ref_clk_clk        => clocks_ref_clk_clk,     --      ref_clk.clk
			ref_reset_reset    => clocks_ref_reset_reset, --    ref_reset.reset
			sys_clk_clk        => clocks_sys_clk_clk,     --      sys_clk.clk
			sdram_clk_clk      => clocks_sdram_clk_clk,   --    sdram_clk.clk
			reset_source_reset => open                    -- reset_source.reset
		);

	cpu : component Nios_System_A1_cpu
		port map (
			clk                                 => clocks_sys_clk_clk,                                --                       clk.clk
			reset_n                             => rst_controller_reset_out_reset_ports_inv,          --                     reset.reset_n
			reset_req                           => rst_controller_reset_out_reset_req,                --                          .reset_req
			d_address                           => cpu_data_master_address,                           --               data_master.address
			d_byteenable                        => cpu_data_master_byteenable,                        --                          .byteenable
			d_read                              => cpu_data_master_read,                              --                          .read
			d_readdata                          => cpu_data_master_readdata,                          --                          .readdata
			d_waitrequest                       => cpu_data_master_waitrequest,                       --                          .waitrequest
			d_write                             => cpu_data_master_write,                             --                          .write
			d_writedata                         => cpu_data_master_writedata,                         --                          .writedata
			debug_mem_slave_debugaccess_to_roms => cpu_data_master_debugaccess,                       --                          .debugaccess
			i_address                           => cpu_instruction_master_address,                    --        instruction_master.address
			i_read                              => cpu_instruction_master_read,                       --                          .read
			i_readdata                          => cpu_instruction_master_readdata,                   --                          .readdata
			i_waitrequest                       => cpu_instruction_master_waitrequest,                --                          .waitrequest
			irq                                 => cpu_irq_irq,                                       --                       irq.irq
			debug_reset_request                 => cpu_debug_reset_request_reset,                     --       debug_reset_request.reset
			debug_mem_slave_address             => mm_interconnect_0_cpu_debug_mem_slave_address,     --           debug_mem_slave.address
			debug_mem_slave_byteenable          => mm_interconnect_0_cpu_debug_mem_slave_byteenable,  --                          .byteenable
			debug_mem_slave_debugaccess         => mm_interconnect_0_cpu_debug_mem_slave_debugaccess, --                          .debugaccess
			debug_mem_slave_read                => mm_interconnect_0_cpu_debug_mem_slave_read,        --                          .read
			debug_mem_slave_readdata            => mm_interconnect_0_cpu_debug_mem_slave_readdata,    --                          .readdata
			debug_mem_slave_waitrequest         => mm_interconnect_0_cpu_debug_mem_slave_waitrequest, --                          .waitrequest
			debug_mem_slave_write               => mm_interconnect_0_cpu_debug_mem_slave_write,       --                          .write
			debug_mem_slave_writedata           => mm_interconnect_0_cpu_debug_mem_slave_writedata,   --                          .writedata
			E_ci_combo_result                   => cpu_custom_instruction_master_result,              -- custom_instruction_master.result
			E_ci_combo_a                        => cpu_custom_instruction_master_a,                   --                          .a
			E_ci_combo_b                        => cpu_custom_instruction_master_b,                   --                          .b
			E_ci_combo_c                        => cpu_custom_instruction_master_c,                   --                          .c
			E_ci_combo_dataa                    => cpu_custom_instruction_master_dataa,               --                          .dataa
			E_ci_combo_datab                    => cpu_custom_instruction_master_datab,               --                          .datab
			E_ci_combo_estatus                  => cpu_custom_instruction_master_estatus,             --                          .estatus
			E_ci_combo_ipending                 => cpu_custom_instruction_master_ipending,            --                          .ipending
			E_ci_combo_n                        => cpu_custom_instruction_master_n,                   --                          .n
			E_ci_combo_readra                   => cpu_custom_instruction_master_readra,              --                          .readra
			E_ci_combo_readrb                   => cpu_custom_instruction_master_readrb,              --                          .readrb
			E_ci_combo_writerc                  => cpu_custom_instruction_master_writerc              --                          .writerc
		);

	high_res_timer : component Nios_System_A1_high_res_timer
		port map (
			clk        => clocks_sys_clk_clk,                                  --   clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,            -- reset.reset_n
			address    => mm_interconnect_0_high_res_timer_s1_address,         --    s1.address
			writedata  => mm_interconnect_0_high_res_timer_s1_writedata,       --      .writedata
			readdata   => mm_interconnect_0_high_res_timer_s1_readdata,        --      .readdata
			chipselect => mm_interconnect_0_high_res_timer_s1_chipselect,      --      .chipselect
			write_n    => mm_interconnect_0_high_res_timer_s1_write_ports_inv, --      .write_n
			irq        => irq_mapper_receiver1_irq                             --   irq.irq
		);

	jtag_uart : component Nios_System_A1_jtag_uart
		port map (
			clk            => clocks_sys_clk_clk,                                            --               clk.clk
			rst_n          => rst_controller_reset_out_reset_ports_inv,                      --             reset.reset_n
			av_chipselect  => mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => mm_interconnect_0_jtag_uart_avalon_jtag_slave_address(0),      --                  .address
			av_read_n      => mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv,  --                  .read_n
			av_readdata    => mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata,        --                  .readdata
			av_write_n     => mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv, --                  .write_n
			av_writedata   => mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata,       --                  .writedata
			av_waitrequest => mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_receiver0_irq                                       --               irq.irq
		);

	onchip_memory : component Nios_System_A1_onchip_memory
		port map (
			clk        => clocks_sys_clk_clk,                            --   clk1.clk
			address    => mm_interconnect_0_onchip_memory_s1_address,    --     s1.address
			clken      => mm_interconnect_0_onchip_memory_s1_clken,      --       .clken
			chipselect => mm_interconnect_0_onchip_memory_s1_chipselect, --       .chipselect
			write      => mm_interconnect_0_onchip_memory_s1_write,      --       .write
			readdata   => mm_interconnect_0_onchip_memory_s1_readdata,   --       .readdata
			writedata  => mm_interconnect_0_onchip_memory_s1_writedata,  --       .writedata
			byteenable => mm_interconnect_0_onchip_memory_s1_byteenable, --       .byteenable
			reset      => rst_controller_reset_out_reset,                -- reset1.reset
			reset_req  => rst_controller_reset_out_reset_req,            --       .reset_req
			freeze     => '0'                                            -- (terminated)
		);

	sdram : component Nios_System_A1_sdram
		port map (
			clk            => clocks_sys_clk_clk,                              --   clk.clk
			reset_n        => rst_controller_reset_out_reset_ports_inv,        -- reset.reset_n
			az_addr        => mm_interconnect_0_sdram_s1_address,              --    s1.address
			az_be_n        => mm_interconnect_0_sdram_s1_byteenable_ports_inv, --      .byteenable_n
			az_cs          => mm_interconnect_0_sdram_s1_chipselect,           --      .chipselect
			az_data        => mm_interconnect_0_sdram_s1_writedata,            --      .writedata
			az_rd_n        => mm_interconnect_0_sdram_s1_read_ports_inv,       --      .read_n
			az_wr_n        => mm_interconnect_0_sdram_s1_write_ports_inv,      --      .write_n
			za_data        => mm_interconnect_0_sdram_s1_readdata,             --      .readdata
			za_valid       => mm_interconnect_0_sdram_s1_readdatavalid,        --      .readdatavalid
			za_waitrequest => mm_interconnect_0_sdram_s1_waitrequest,          --      .waitrequest
			zs_addr        => sdram_wire_addr,                                 --  wire.export
			zs_ba          => sdram_wire_ba,                                   --      .export
			zs_cas_n       => sdram_wire_cas_n,                                --      .export
			zs_cke         => sdram_wire_cke,                                  --      .export
			zs_cs_n        => sdram_wire_cs_n,                                 --      .export
			zs_dq          => sdram_wire_dq,                                   --      .export
			zs_dqm         => sdram_wire_dqm,                                  --      .export
			zs_ras_n       => sdram_wire_ras_n,                                --      .export
			zs_we_n        => sdram_wire_we_n                                  --      .export
		);

	cpu_custom_instruction_master_translator : component altera_customins_master_translator
		generic map (
			SHARED_COMB_AND_MULTI => 0
		)
		port map (
			ci_slave_dataa            => cpu_custom_instruction_master_dataa,                              --       ci_slave.dataa
			ci_slave_datab            => cpu_custom_instruction_master_datab,                              --               .datab
			ci_slave_result           => cpu_custom_instruction_master_result,                             --               .result
			ci_slave_n                => cpu_custom_instruction_master_n,                                  --               .n
			ci_slave_readra           => cpu_custom_instruction_master_readra,                             --               .readra
			ci_slave_readrb           => cpu_custom_instruction_master_readrb,                             --               .readrb
			ci_slave_writerc          => cpu_custom_instruction_master_writerc,                            --               .writerc
			ci_slave_a                => cpu_custom_instruction_master_a,                                  --               .a
			ci_slave_b                => cpu_custom_instruction_master_b,                                  --               .b
			ci_slave_c                => cpu_custom_instruction_master_c,                                  --               .c
			ci_slave_ipending         => cpu_custom_instruction_master_ipending,                           --               .ipending
			ci_slave_estatus          => cpu_custom_instruction_master_estatus,                            --               .estatus
			comb_ci_master_dataa      => cpu_custom_instruction_master_translator_comb_ci_master_dataa,    -- comb_ci_master.dataa
			comb_ci_master_datab      => cpu_custom_instruction_master_translator_comb_ci_master_datab,    --               .datab
			comb_ci_master_result     => cpu_custom_instruction_master_translator_comb_ci_master_result,   --               .result
			comb_ci_master_n          => cpu_custom_instruction_master_translator_comb_ci_master_n,        --               .n
			comb_ci_master_readra     => cpu_custom_instruction_master_translator_comb_ci_master_readra,   --               .readra
			comb_ci_master_readrb     => cpu_custom_instruction_master_translator_comb_ci_master_readrb,   --               .readrb
			comb_ci_master_writerc    => cpu_custom_instruction_master_translator_comb_ci_master_writerc,  --               .writerc
			comb_ci_master_a          => cpu_custom_instruction_master_translator_comb_ci_master_a,        --               .a
			comb_ci_master_b          => cpu_custom_instruction_master_translator_comb_ci_master_b,        --               .b
			comb_ci_master_c          => cpu_custom_instruction_master_translator_comb_ci_master_c,        --               .c
			comb_ci_master_ipending   => cpu_custom_instruction_master_translator_comb_ci_master_ipending, --               .ipending
			comb_ci_master_estatus    => cpu_custom_instruction_master_translator_comb_ci_master_estatus,  --               .estatus
			ci_slave_multi_clk        => '0',                                                              --    (terminated)
			ci_slave_multi_reset      => '0',                                                              --    (terminated)
			ci_slave_multi_clken      => '0',                                                              --    (terminated)
			ci_slave_multi_reset_req  => '0',                                                              --    (terminated)
			ci_slave_multi_start      => '0',                                                              --    (terminated)
			ci_slave_multi_done       => open,                                                             --    (terminated)
			ci_slave_multi_dataa      => "00000000000000000000000000000000",                               --    (terminated)
			ci_slave_multi_datab      => "00000000000000000000000000000000",                               --    (terminated)
			ci_slave_multi_result     => open,                                                             --    (terminated)
			ci_slave_multi_n          => "00000000",                                                       --    (terminated)
			ci_slave_multi_readra     => '0',                                                              --    (terminated)
			ci_slave_multi_readrb     => '0',                                                              --    (terminated)
			ci_slave_multi_writerc    => '0',                                                              --    (terminated)
			ci_slave_multi_a          => "00000",                                                          --    (terminated)
			ci_slave_multi_b          => "00000",                                                          --    (terminated)
			ci_slave_multi_c          => "00000",                                                          --    (terminated)
			multi_ci_master_clk       => open,                                                             --    (terminated)
			multi_ci_master_reset     => open,                                                             --    (terminated)
			multi_ci_master_clken     => open,                                                             --    (terminated)
			multi_ci_master_reset_req => open,                                                             --    (terminated)
			multi_ci_master_start     => open,                                                             --    (terminated)
			multi_ci_master_done      => '0',                                                              --    (terminated)
			multi_ci_master_dataa     => open,                                                             --    (terminated)
			multi_ci_master_datab     => open,                                                             --    (terminated)
			multi_ci_master_result    => "00000000000000000000000000000000",                               --    (terminated)
			multi_ci_master_n         => open,                                                             --    (terminated)
			multi_ci_master_readra    => open,                                                             --    (terminated)
			multi_ci_master_readrb    => open,                                                             --    (terminated)
			multi_ci_master_writerc   => open,                                                             --    (terminated)
			multi_ci_master_a         => open,                                                             --    (terminated)
			multi_ci_master_b         => open,                                                             --    (terminated)
			multi_ci_master_c         => open                                                              --    (terminated)
		);

	cpu_custom_instruction_master_comb_xconnect : component Nios_System_A1_cpu_custom_instruction_master_comb_xconnect
		port map (
			ci_slave_dataa      => cpu_custom_instruction_master_translator_comb_ci_master_dataa,    --   ci_slave.dataa
			ci_slave_datab      => cpu_custom_instruction_master_translator_comb_ci_master_datab,    --           .datab
			ci_slave_result     => cpu_custom_instruction_master_translator_comb_ci_master_result,   --           .result
			ci_slave_n          => cpu_custom_instruction_master_translator_comb_ci_master_n,        --           .n
			ci_slave_readra     => cpu_custom_instruction_master_translator_comb_ci_master_readra,   --           .readra
			ci_slave_readrb     => cpu_custom_instruction_master_translator_comb_ci_master_readrb,   --           .readrb
			ci_slave_writerc    => cpu_custom_instruction_master_translator_comb_ci_master_writerc,  --           .writerc
			ci_slave_a          => cpu_custom_instruction_master_translator_comb_ci_master_a,        --           .a
			ci_slave_b          => cpu_custom_instruction_master_translator_comb_ci_master_b,        --           .b
			ci_slave_c          => cpu_custom_instruction_master_translator_comb_ci_master_c,        --           .c
			ci_slave_ipending   => cpu_custom_instruction_master_translator_comb_ci_master_ipending, --           .ipending
			ci_slave_estatus    => cpu_custom_instruction_master_translator_comb_ci_master_estatus,  --           .estatus
			ci_master0_dataa    => cpu_custom_instruction_master_comb_xconnect_ci_master0_dataa,     -- ci_master0.dataa
			ci_master0_datab    => cpu_custom_instruction_master_comb_xconnect_ci_master0_datab,     --           .datab
			ci_master0_result   => cpu_custom_instruction_master_comb_xconnect_ci_master0_result,    --           .result
			ci_master0_n        => cpu_custom_instruction_master_comb_xconnect_ci_master0_n,         --           .n
			ci_master0_readra   => cpu_custom_instruction_master_comb_xconnect_ci_master0_readra,    --           .readra
			ci_master0_readrb   => cpu_custom_instruction_master_comb_xconnect_ci_master0_readrb,    --           .readrb
			ci_master0_writerc  => cpu_custom_instruction_master_comb_xconnect_ci_master0_writerc,   --           .writerc
			ci_master0_a        => cpu_custom_instruction_master_comb_xconnect_ci_master0_a,         --           .a
			ci_master0_b        => cpu_custom_instruction_master_comb_xconnect_ci_master0_b,         --           .b
			ci_master0_c        => cpu_custom_instruction_master_comb_xconnect_ci_master0_c,         --           .c
			ci_master0_ipending => cpu_custom_instruction_master_comb_xconnect_ci_master0_ipending,  --           .ipending
			ci_master0_estatus  => cpu_custom_instruction_master_comb_xconnect_ci_master0_estatus    --           .estatus
		);

	cpu_custom_instruction_master_comb_slave_translator0 : component altera_customins_slave_translator
		generic map (
			N_WIDTH          => 8,
			USE_DONE         => 0,
			NUM_FIXED_CYCLES => 0
		)
		port map (
			ci_slave_dataa      => cpu_custom_instruction_master_comb_xconnect_ci_master0_dataa,          --  ci_slave.dataa
			ci_slave_datab      => cpu_custom_instruction_master_comb_xconnect_ci_master0_datab,          --          .datab
			ci_slave_result     => cpu_custom_instruction_master_comb_xconnect_ci_master0_result,         --          .result
			ci_slave_n          => cpu_custom_instruction_master_comb_xconnect_ci_master0_n,              --          .n
			ci_slave_readra     => cpu_custom_instruction_master_comb_xconnect_ci_master0_readra,         --          .readra
			ci_slave_readrb     => cpu_custom_instruction_master_comb_xconnect_ci_master0_readrb,         --          .readrb
			ci_slave_writerc    => cpu_custom_instruction_master_comb_xconnect_ci_master0_writerc,        --          .writerc
			ci_slave_a          => cpu_custom_instruction_master_comb_xconnect_ci_master0_a,              --          .a
			ci_slave_b          => cpu_custom_instruction_master_comb_xconnect_ci_master0_b,              --          .b
			ci_slave_c          => cpu_custom_instruction_master_comb_xconnect_ci_master0_c,              --          .c
			ci_slave_ipending   => cpu_custom_instruction_master_comb_xconnect_ci_master0_ipending,       --          .ipending
			ci_slave_estatus    => cpu_custom_instruction_master_comb_xconnect_ci_master0_estatus,        --          .estatus
			ci_master_dataa     => cpu_custom_instruction_master_comb_slave_translator0_ci_master_dataa,  -- ci_master.dataa
			ci_master_datab     => cpu_custom_instruction_master_comb_slave_translator0_ci_master_datab,  --          .datab
			ci_master_result    => cpu_custom_instruction_master_comb_slave_translator0_ci_master_result, --          .result
			ci_master_n         => open,                                                                  -- (terminated)
			ci_master_readra    => open,                                                                  -- (terminated)
			ci_master_readrb    => open,                                                                  -- (terminated)
			ci_master_writerc   => open,                                                                  -- (terminated)
			ci_master_a         => open,                                                                  -- (terminated)
			ci_master_b         => open,                                                                  -- (terminated)
			ci_master_c         => open,                                                                  -- (terminated)
			ci_master_ipending  => open,                                                                  -- (terminated)
			ci_master_estatus   => open,                                                                  -- (terminated)
			ci_master_clk       => open,                                                                  -- (terminated)
			ci_master_clken     => open,                                                                  -- (terminated)
			ci_master_reset_req => open,                                                                  -- (terminated)
			ci_master_reset     => open,                                                                  -- (terminated)
			ci_master_start     => open,                                                                  -- (terminated)
			ci_master_done      => '0',                                                                   -- (terminated)
			ci_slave_clk        => '0',                                                                   -- (terminated)
			ci_slave_clken      => '0',                                                                   -- (terminated)
			ci_slave_reset_req  => '0',                                                                   -- (terminated)
			ci_slave_reset      => '0',                                                                   -- (terminated)
			ci_slave_start      => '0',                                                                   -- (terminated)
			ci_slave_done       => open                                                                   -- (terminated)
		);

	mm_interconnect_0 : component Nios_System_A1_mm_interconnect_0
		port map (
			clocks_sys_clk_clk                      => clocks_sys_clk_clk,                                        --                  clocks_sys_clk.clk
			cpu_reset_reset_bridge_in_reset_reset   => rst_controller_reset_out_reset,                            -- cpu_reset_reset_bridge_in_reset.reset
			cpu_data_master_address                 => cpu_data_master_address,                                   --                 cpu_data_master.address
			cpu_data_master_waitrequest             => cpu_data_master_waitrequest,                               --                                .waitrequest
			cpu_data_master_byteenable              => cpu_data_master_byteenable,                                --                                .byteenable
			cpu_data_master_read                    => cpu_data_master_read,                                      --                                .read
			cpu_data_master_readdata                => cpu_data_master_readdata,                                  --                                .readdata
			cpu_data_master_write                   => cpu_data_master_write,                                     --                                .write
			cpu_data_master_writedata               => cpu_data_master_writedata,                                 --                                .writedata
			cpu_data_master_debugaccess             => cpu_data_master_debugaccess,                               --                                .debugaccess
			cpu_instruction_master_address          => cpu_instruction_master_address,                            --          cpu_instruction_master.address
			cpu_instruction_master_waitrequest      => cpu_instruction_master_waitrequest,                        --                                .waitrequest
			cpu_instruction_master_read             => cpu_instruction_master_read,                               --                                .read
			cpu_instruction_master_readdata         => cpu_instruction_master_readdata,                           --                                .readdata
			BUTTON_pio_s1_address                   => mm_interconnect_0_button_pio_s1_address,                   --                   BUTTON_pio_s1.address
			BUTTON_pio_s1_write                     => mm_interconnect_0_button_pio_s1_write,                     --                                .write
			BUTTON_pio_s1_readdata                  => mm_interconnect_0_button_pio_s1_readdata,                  --                                .readdata
			BUTTON_pio_s1_writedata                 => mm_interconnect_0_button_pio_s1_writedata,                 --                                .writedata
			BUTTON_pio_s1_chipselect                => mm_interconnect_0_button_pio_s1_chipselect,                --                                .chipselect
			cpu_debug_mem_slave_address             => mm_interconnect_0_cpu_debug_mem_slave_address,             --             cpu_debug_mem_slave.address
			cpu_debug_mem_slave_write               => mm_interconnect_0_cpu_debug_mem_slave_write,               --                                .write
			cpu_debug_mem_slave_read                => mm_interconnect_0_cpu_debug_mem_slave_read,                --                                .read
			cpu_debug_mem_slave_readdata            => mm_interconnect_0_cpu_debug_mem_slave_readdata,            --                                .readdata
			cpu_debug_mem_slave_writedata           => mm_interconnect_0_cpu_debug_mem_slave_writedata,           --                                .writedata
			cpu_debug_mem_slave_byteenable          => mm_interconnect_0_cpu_debug_mem_slave_byteenable,          --                                .byteenable
			cpu_debug_mem_slave_waitrequest         => mm_interconnect_0_cpu_debug_mem_slave_waitrequest,         --                                .waitrequest
			cpu_debug_mem_slave_debugaccess         => mm_interconnect_0_cpu_debug_mem_slave_debugaccess,         --                                .debugaccess
			high_res_timer_s1_address               => mm_interconnect_0_high_res_timer_s1_address,               --               high_res_timer_s1.address
			high_res_timer_s1_write                 => mm_interconnect_0_high_res_timer_s1_write,                 --                                .write
			high_res_timer_s1_readdata              => mm_interconnect_0_high_res_timer_s1_readdata,              --                                .readdata
			high_res_timer_s1_writedata             => mm_interconnect_0_high_res_timer_s1_writedata,             --                                .writedata
			high_res_timer_s1_chipselect            => mm_interconnect_0_high_res_timer_s1_chipselect,            --                                .chipselect
			jtag_uart_avalon_jtag_slave_address     => mm_interconnect_0_jtag_uart_avalon_jtag_slave_address,     --     jtag_uart_avalon_jtag_slave.address
			jtag_uart_avalon_jtag_slave_write       => mm_interconnect_0_jtag_uart_avalon_jtag_slave_write,       --                                .write
			jtag_uart_avalon_jtag_slave_read        => mm_interconnect_0_jtag_uart_avalon_jtag_slave_read,        --                                .read
			jtag_uart_avalon_jtag_slave_readdata    => mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata,    --                                .readdata
			jtag_uart_avalon_jtag_slave_writedata   => mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata,   --                                .writedata
			jtag_uart_avalon_jtag_slave_waitrequest => mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest, --                                .waitrequest
			jtag_uart_avalon_jtag_slave_chipselect  => mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect,  --                                .chipselect
			LED_pio_s1_address                      => mm_interconnect_0_led_pio_s1_address,                      --                      LED_pio_s1.address
			LED_pio_s1_write                        => mm_interconnect_0_led_pio_s1_write,                        --                                .write
			LED_pio_s1_readdata                     => mm_interconnect_0_led_pio_s1_readdata,                     --                                .readdata
			LED_pio_s1_writedata                    => mm_interconnect_0_led_pio_s1_writedata,                    --                                .writedata
			LED_pio_s1_chipselect                   => mm_interconnect_0_led_pio_s1_chipselect,                   --                                .chipselect
			onchip_memory_s1_address                => mm_interconnect_0_onchip_memory_s1_address,                --                onchip_memory_s1.address
			onchip_memory_s1_write                  => mm_interconnect_0_onchip_memory_s1_write,                  --                                .write
			onchip_memory_s1_readdata               => mm_interconnect_0_onchip_memory_s1_readdata,               --                                .readdata
			onchip_memory_s1_writedata              => mm_interconnect_0_onchip_memory_s1_writedata,              --                                .writedata
			onchip_memory_s1_byteenable             => mm_interconnect_0_onchip_memory_s1_byteenable,             --                                .byteenable
			onchip_memory_s1_chipselect             => mm_interconnect_0_onchip_memory_s1_chipselect,             --                                .chipselect
			onchip_memory_s1_clken                  => mm_interconnect_0_onchip_memory_s1_clken,                  --                                .clken
			sdram_s1_address                        => mm_interconnect_0_sdram_s1_address,                        --                        sdram_s1.address
			sdram_s1_write                          => mm_interconnect_0_sdram_s1_write,                          --                                .write
			sdram_s1_read                           => mm_interconnect_0_sdram_s1_read,                           --                                .read
			sdram_s1_readdata                       => mm_interconnect_0_sdram_s1_readdata,                       --                                .readdata
			sdram_s1_writedata                      => mm_interconnect_0_sdram_s1_writedata,                      --                                .writedata
			sdram_s1_byteenable                     => mm_interconnect_0_sdram_s1_byteenable,                     --                                .byteenable
			sdram_s1_readdatavalid                  => mm_interconnect_0_sdram_s1_readdatavalid,                  --                                .readdatavalid
			sdram_s1_waitrequest                    => mm_interconnect_0_sdram_s1_waitrequest,                    --                                .waitrequest
			sdram_s1_chipselect                     => mm_interconnect_0_sdram_s1_chipselect,                     --                                .chipselect
			Segment_1_s1_address                    => mm_interconnect_0_segment_1_s1_address,                    --                    Segment_1_s1.address
			Segment_1_s1_write                      => mm_interconnect_0_segment_1_s1_write,                      --                                .write
			Segment_1_s1_readdata                   => mm_interconnect_0_segment_1_s1_readdata,                   --                                .readdata
			Segment_1_s1_writedata                  => mm_interconnect_0_segment_1_s1_writedata,                  --                                .writedata
			Segment_1_s1_chipselect                 => mm_interconnect_0_segment_1_s1_chipselect,                 --                                .chipselect
			Segment_2_s1_address                    => mm_interconnect_0_segment_2_s1_address,                    --                    Segment_2_s1.address
			Segment_2_s1_write                      => mm_interconnect_0_segment_2_s1_write,                      --                                .write
			Segment_2_s1_readdata                   => mm_interconnect_0_segment_2_s1_readdata,                   --                                .readdata
			Segment_2_s1_writedata                  => mm_interconnect_0_segment_2_s1_writedata,                  --                                .writedata
			Segment_2_s1_chipselect                 => mm_interconnect_0_segment_2_s1_chipselect,                 --                                .chipselect
			Segment_3_s1_address                    => mm_interconnect_0_segment_3_s1_address,                    --                    Segment_3_s1.address
			Segment_3_s1_write                      => mm_interconnect_0_segment_3_s1_write,                      --                                .write
			Segment_3_s1_readdata                   => mm_interconnect_0_segment_3_s1_readdata,                   --                                .readdata
			Segment_3_s1_writedata                  => mm_interconnect_0_segment_3_s1_writedata,                  --                                .writedata
			Segment_3_s1_chipselect                 => mm_interconnect_0_segment_3_s1_chipselect,                 --                                .chipselect
			Segment_4_s1_address                    => mm_interconnect_0_segment_4_s1_address,                    --                    Segment_4_s1.address
			Segment_4_s1_write                      => mm_interconnect_0_segment_4_s1_write,                      --                                .write
			Segment_4_s1_readdata                   => mm_interconnect_0_segment_4_s1_readdata,                   --                                .readdata
			Segment_4_s1_writedata                  => mm_interconnect_0_segment_4_s1_writedata,                  --                                .writedata
			Segment_4_s1_chipselect                 => mm_interconnect_0_segment_4_s1_chipselect,                 --                                .chipselect
			Switches_0_7_s1_address                 => mm_interconnect_0_switches_0_7_s1_address,                 --                 Switches_0_7_s1.address
			Switches_0_7_s1_readdata                => mm_interconnect_0_switches_0_7_s1_readdata                 --                                .readdata
		);

	irq_mapper : component Nios_System_A1_irq_mapper
		port map (
			clk           => clocks_sys_clk_clk,             --       clk.clk
			reset         => rst_controller_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,       -- receiver0.irq
			receiver1_irq => irq_mapper_receiver1_irq,       -- receiver1.irq
			receiver2_irq => irq_mapper_receiver2_irq,       -- receiver2.irq
			sender_irq    => cpu_irq_irq                     --    sender.irq
		);

	rst_controller : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => cpu_debug_reset_request_reset,      -- reset_in0.reset
			clk            => clocks_sys_clk_clk,                 --       clk.clk
			reset_out      => rst_controller_reset_out_reset,     -- reset_out.reset
			reset_req      => rst_controller_reset_out_reset_req, --          .reset_req
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv <= not mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;

	mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv <= not mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;

	mm_interconnect_0_led_pio_s1_write_ports_inv <= not mm_interconnect_0_led_pio_s1_write;

	mm_interconnect_0_sdram_s1_read_ports_inv <= not mm_interconnect_0_sdram_s1_read;

	mm_interconnect_0_sdram_s1_byteenable_ports_inv <= not mm_interconnect_0_sdram_s1_byteenable;

	mm_interconnect_0_sdram_s1_write_ports_inv <= not mm_interconnect_0_sdram_s1_write;

	mm_interconnect_0_high_res_timer_s1_write_ports_inv <= not mm_interconnect_0_high_res_timer_s1_write;

	mm_interconnect_0_button_pio_s1_write_ports_inv <= not mm_interconnect_0_button_pio_s1_write;

	mm_interconnect_0_segment_1_s1_write_ports_inv <= not mm_interconnect_0_segment_1_s1_write;

	mm_interconnect_0_segment_2_s1_write_ports_inv <= not mm_interconnect_0_segment_2_s1_write;

	mm_interconnect_0_segment_3_s1_write_ports_inv <= not mm_interconnect_0_segment_3_s1_write;

	mm_interconnect_0_segment_4_s1_write_ports_inv <= not mm_interconnect_0_segment_4_s1_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

end architecture rtl; -- of Nios_System_A1
